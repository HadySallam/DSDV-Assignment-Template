module template_tb;
  logic a, b, c, d, e;
  logic z;

  template DUT (.a(a), .b(b), .c(c), .d(d), .e(e), .z(z));

  initial
    begin

    end
endmodule
