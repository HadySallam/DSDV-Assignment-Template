module template(input a, b, c, d, e
                output z);
  
end module
